module bin_bindec(
	input 	[5:0]	bin,
	output	[3:0]	bindec_first,
	output	[3:0]	bindec_second
);

	


endmodule;