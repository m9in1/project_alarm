`define APB_WIDTH 32
`define DIS_FREQ 22000


module sound(
	input clk,
	input [`APB_WIDTH-1:0] 	datadig_i,
	output [`APB_WIDTH-1:0]	dataan_o,
	output data_ready
	);

	
endmodule;